module io();
  //inout [7:0] databus;
  //output ior, iow;
  //reg [7:0] idr;
endmodule
